`include "full_substractor.v"


module full_subtractor_64_bit();
endmodule