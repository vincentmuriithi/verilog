module dFlipFlop(A,D, CLK);
endmodule
