`include "full_subtractor.v"


module full_subtractor_64_bit();
endmodule