module gate1;
endmodule